// $Id: $
// File name:   mealy.sv
// Created:     2/9/2016
// Author:      Arnav Mittal
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: This is the mealy diagram
