// Description: This is the test bench for the Slave Inner block
`timescale 1ns / 10ps

module tb_slave_inner();
  
  // Define parameters
	parameter CLK_PERIOD	= 10;
	parameter SCL_PERIOD    = 300;
	parameter sclwait       = 300;
  
	reg tb_clk;
  reg tb_n_rst;
  reg [7:0] tb_tx_data;   // Data coming in from the TX FIFO
  reg tb_address_mode;
  reg tb_ms_select;
  reg [9:0] tb_bus_address;
  reg tb_en_clock_strech;
  reg tb_TX_fifo_empty;
  reg tb_RX_fifo_full;
  reg tb_RX_fifo_almost_full;
  reg tb_SDA_sync;
  reg tb_SCL_sync;
  reg [7:0] tb_rx_data_slave;
  reg tb_set_transaction_complete_slave;
  reg tb_ack_error_set_slave;
  reg tb_busy_slave;
  reg tb_TX_read_enable_slave;
  reg tb_RX_write_enable_slave;
  reg tb_SDA_out_slave;
  reg tb_SCL_sync_out_slave;

	slave_inner SLAVE_INNER
	(
		.clk(tb_clk),
    .n_rst(tb_n_rst),
    .tx_data(tb_tx_data),
    .address_mode(tb_address_mode),
    .ms_select(tb_ms_select),
    .bus_address(tb_bus_address),
    .en_clock_strech(tb_en_clock_strech),
    .TX_fifo_empty(tb_TX_fifo_empty),
    .RX_fifo_full(tb_RX_fifo_full),
    .RX_fifo_almost_full(tb_RX_fifo_almost_full),
    .SDA_sync(tb_SDA_sync),
    .SCL_sync(tb_SCL_sync),
    .rx_data_slave(tb_rx_data_slave),
    .set_transaction_complete_slave(tb_set_transaction_complete_slave),
    .ack_error_set_slave(tb_ack_error_set_slave),
    .busy_slave(tb_busy_slave),
    .TX_read_enable_slave(tb_TX_read_enable_slave),
    .RX_write_enable_slave(tb_RX_write_enable_slave),
    .SDA_out_slave(tb_SDA_out_slave),
    .SCL_out_slave(tb_SCL_sync_out_slave)
	);
	
	always
	begin : CLK_GEN
		tb_clk = 1'b0;
		#(CLK_PERIOD / 2);
		tb_clk = 1'b1;
		#(CLK_PERIOD / 2);
	end
	
	always
	begin : SCL_GEN
	    tb_SCL_sync = 1'b0;
	    #(SCL_PERIOD / 3);
	    tb_SCL_sync = 1'b1;
	    #(SCL_PERIOD / 3); 
	    tb_SCL_sync = 1'b0;
	    #(SCL_PERIOD / 3);
	end	
  
  integer i;

	initial
	begin 
	  tb_n_rst = 1'b0;
    tb_tx_data = 8'b00000000;
    tb_address_mode = 1'b0;   // 7 Bit Mode 
    tb_ms_select = 1'b0;      // Slave selected
    tb_bus_address = 10'b0000000111;
    tb_en_clock_strech = 1'b0;
    tb_TX_fifo_empty = 1'b0;
    tb_RX_fifo_full = 1'b0;
    tb_RX_fifo_almost_full = 1'b0;
    tb_SDA_sync = 1'b0;
	  @(posedge tb_clk);
    tb_n_rst = 1'b1;
 
    
    @(posedge tb_clk);
    @(posedge tb_clk);
    @(posedge tb_clk);
    @(posedge tb_clk);
    @(posedge tb_clk); 
    
    // Generate a Start Condition by varying SDA line.
    tb_SDA_sync = 1'b1;

    @(posedge tb_SCL_sync);
    @(posedge tb_clk);
    @(posedge tb_clk);
    @(posedge tb_clk);
    @(posedge tb_clk);
    @(posedge tb_clk);

    tb_SDA_sync = 1'b0;

    i=0;
    repeat (20) 
    begin
      @(negedge tb_SCL_sync);
      i = i+1;
      tb_SDA_sync = 1'b0;
      if(i == 19) 
      begin
         @(posedge tb_SCL_sync);
         @(posedge tb_clk);
         @(posedge tb_clk);
         tb_SDA_sync = 1'b1;
       end 
    end

    // Set bus_address = 0001100110.
    // Send address 7 bit '1100110'+'1' denoting read from SDA line.
    // Check if Ack sent by slave on 9th pulse of SCL line.
    
    
	end 
endmodule
