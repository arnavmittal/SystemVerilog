/home/ecegrid/a/mg150/ece337/Lab2/source/tb_adder_nbit.sv