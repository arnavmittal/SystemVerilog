// $Id: $
// File name:   shift_register.sv
// Created:     2/26/2016
// Author:      Arnav Mittal
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: This is the module for the Shift register of the USB Receiver Lab
//              which hold the 1 byte of data to be stored in the FIFO.
