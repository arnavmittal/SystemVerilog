/home/ecegrid/a/mg150/ece337/Lab2/source/adder_8bit.sv